package spi_env_pkg;
  import uvm_pkg::*;
  `include "uvm_macros.svh"

  import spi_common_agent_pkg::*;
  import spi_m_agent_pkg::*;
  import spi_ms_agent_pkg::*;
  `include "spi_env.sv"
endpackage