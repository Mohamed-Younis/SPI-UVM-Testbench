package spi_env_pkg;
  import uvm_pkg::*;
  `include "uvm_macros.svh"

  import spi_common_agent_pkg::*;
  import spi_s_agent_pkg::*;
  import spi_sm_agent_pkg::*;
  `include "spi_scoreboard.sv"
  `include "spi_env.sv"
endpackage