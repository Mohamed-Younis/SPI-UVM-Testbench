package spi_common_agent_pkg;
  import uvm_pkg::*;
  `include "uvm_macros.svh"

  `include "spi_seq_item.sv"
  `include "spi_sequence.sv"
endpackage