package master_slave_spi_test_pkg;
  import uvm_pkg::*;
  `include "uvm_macros.svh"

  import spi_common_agent_pkg::*;
  import spi_m_agent_pkg::*;
  import spi_s_agent_pkg::*;
  import spi_ms_agent_pkg::*;
  import master_slave_spi_env_pkg::*;

  `include "master_slave_spi_base_test.sv"
endpackage