package spi_test_pkg;
  import uvm_pkg::*;
  `include "uvm_macros.svh"

  import spi_common_agent_pkg::*;
  import spi_s_agent_pkg::*;
  import spi_sm_agent_pkg::*;
  import spi_env_pkg::*;

  `include "spi_base_test.sv"
endpackage